module transcodor (input [6:0] s,
						 output reg [13:0] q);
	
			always@(s)
				case(s)
					  0: q=14'b10000001000000;
					  1: q=14'b10000001111001;
					  2: q=14'b10000000100100;
					  3: q=14'b10000000110000;
					  4: q=14'b10000000011001;
					  5: q=14'b10000000010010;
					  6: q=14'b10000000000010;
					  7: q=14'b10000001111000;
					  8: q=14'b10000000000000;
					  9: q=14'b10000000010000;
					  10: q=14'b11110011000000;
					  11: q=14'b11110011111001;
					  12: q=14'b11110010100100;
					  13: q=14'b11110010110000;
					  14: q=14'b11110010011001;
					  15: q=14'b11110010010010;
					  16: q=14'b11110010000010;
					  17: q=14'b11110011111000;
					  18: q=14'b11110010000000;
					  19: q=14'b11110010010000;
					  20: q=14'b01001001000000;
					  21: q=14'b01001001111001;
					  22: q=14'b01001000100100;
					  23: q=14'b01001000110000;
					  24: q=14'b01001000011001;
					  25: q=14'b01001000010010;
					  26: q=14'b01001000000010;
					  27: q=14'b01001001111000;
					  28: q=14'b01001000000000;
					  29: q=14'b01001000010000;
					  30: q=14'b01100001000000;
					  31: q=14'b01100001111001;
					  32: q=14'b01100000100100;
					  33: q=14'b01100000110000;
					  34: q=14'b01100000011001;
					  35: q=14'b01100000010010;
					  36: q=14'b01100000000010;
					  37: q=14'b01100001111000;
					  38: q=14'b01100000000000;
					  39: q=14'b01100000010000;
					  40: q=14'b00110011000000;
					  41: q=14'b00110011111001;
					  42: q=14'b00110010100100;
					  43: q=14'b00110010110000;
					  44: q=14'b00110010011001;
					  45: q=14'b00110010010010;
					  46: q=14'b00110010000010;
					  47: q=14'b00110011111000;
					  48: q=14'b00110010000000;
					  49: q=14'b00110010010000;
					  50: q=14'b00100101000000;
					  51: q=14'b00100101111001;
					  52: q=14'b00100100100100;
					  53: q=14'b00100100110000;
					  54: q=14'b00100100011001;
					  55: q=14'b00100100010010;
					  56: q=14'b00100100000010;
					  57: q=14'b00100101111000;
					  58: q=14'b00100100000000;
					  59: q=14'b00100100010000;
					  60: q=14'b00000101000000;
					  61: q=14'b00000101111001;
					  62: q=14'b00000100100100;
					  63: q=14'b00000100110000;
					  
					  default:
					  q=14'b10000001111001;
					  
				endcase
			
endmodule